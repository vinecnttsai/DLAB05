/*
  BCD_seq: Sequential BCD Display Controller
  ------------------------------------------

  Description:
    This top-level module integrates a 4-bit up/down counter, a frequency divider,
    and a 7-segment decoder to control a BCD output display.
    It uses a slow clock (1 Hz) generated from the 100 MHz input clock to drive
    the counter, and then decodes the counter output to display it on a 7-segment display.

  Modules Used:
    - fq_div: Frequency divider that converts 100 MHz input clock to 1 Hz
    - cnt_4b: 4-bit up/down counter (parameterized with Max=15, Min=0)
    - svn_dcdr: 7-segment decoder with digit selection and decimal point control

  Ports:
    Inputs:
      - clk100M   : 100 MHz system clock
      - sys_rst_n : Active-low asynchronous reset
      - dp_in     : Decimal point control input
      - U_D       : Count direction control (1 = up, 0 = down)
    Outputs:
      - CA to CG  : Segment outputs (7-segment display)
      - DP        : Decimal point output
      - AN[7:0]   : Digit enable outputs (for multiplexed displays)

  Internal Signals:
    - clk  : 1 Hz clock generated by fq_div
    - cnt  : 4-bit counter output (0~15)

*/

module BCD_seq (
    input clk100M,
    input sys_rst_n,
    input dp_in,
    input U_D,
    output CA, 
    output CB,
    output CC, 
    output CD, 
    output CE,
    output CF, 
    output CG,
    output DP,
    output [7:0] AN
);
wire clk;
wire [3:0] cnt;

(* keep_hierarchy = "yes" *)svn_dcdr svn1 (
    .in(cnt),
    .dp_in(dp_in),
    .CA(CA),
    .CB(CB),
    .CC(CC),
    .CD(CD),
    .CE(CE),
    .CF(CF),
    .CG(CG),
    .DP(DP),
    .AN(AN)
);

(* keep_hierarchy = "yes" *)fq_div #(100_000_000) fq_div_100M (
    .rst_n(sys_rst_n),
    .org_clk(clk100M),
    .div_n_clk(clk)
);

(* keep_hierarchy = "yes" *)cnt_4b #(.Max(15), .Min(0)) cnt_9 (
    .clk(clk),
    .rst_n(sys_rst_n),
    .U_D(U_D),
    .cnt(cnt)
);
assign out = cnt;

endmodule
